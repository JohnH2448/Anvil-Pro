package Configuration;

    parameter [31:0] resetVector = 32'd0;

endpackage
