typedef struct packed {
    logic [3:0] ageTag;
    logic isLoad;
    logic busy;
} RegisterStatusEntry_;